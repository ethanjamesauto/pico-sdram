`timescale 1ns / 1ps

module test_sdram;

/*
module MT48LC8M16A2 (dq, addr, ba, clk, cke, csb, rasb, casb, web, dqm);

    parameter addr_bits =      13;
    parameter data_bits =      16;
    parameter col_bits  =       9;
    parameter mem_sizes = 2097151;                                  // 2 Meg
 
    inout     [data_bits - 1 : 0] dq;
    input     [addr_bits - 1 : 0] addr;
    input                 [1 : 0] ba;
    input                         clk;
    input                         cke;
    input                         csb;
    input                         rasb;
    input                         casb;
    input                         web;
    input                 [1 : 0] dqm;
*/

wire [15:0] dq;
logic [12:0] addr;
logic [1:0] ba;
logic clk;
logic cke;
logic csb;
logic rasb;
logic casb;
logic web;
logic [1:0] dqm;

logic srclk, rclk, ser1, ser2, ser3;

assign srclk = clk;
assign csb = rclk;

IS42VM16400K
// MT48LC8M16A2 
sdram(
    .dq(dq),
    .addr(addr),
    .ba(ba),
    .clk(clk),
    .cke(cke),
    .csb(csb),
    .rasb(rasb),
    .casb(casb),
    .web(web),
    .dqm(dqm)
);

\74595 one(
    .SER(ser1),
    .SCLK(srclk),
    .RCLK(rclk),
    .OE_n(1'b0),
    .CLR_n(1'b1),
    .VCC(1'b1),
    .GND(1'b0),
    .Q_A(addr[4]),
    .Q_B(addr[12]),
    .Q_C(addr[11]),
    .Q_D(addr[9]),
    .Q_E(addr[8]),
    .Q_F(addr[7]),
    .Q_G(addr[6]),
    .Q_H(addr[5]),
    .Q_H_n()
);

\74595 two(
    .SER(ser2),
    .SCLK(srclk),
    .RCLK(rclk),
    .OE_n(1'b0),
    .CLR_n(1'b1),
    .VCC(1'b1),
    .GND(1'b0),
    .Q_A(ba[0]),
    .Q_B(),
    .Q_C(addr[3]),
    .Q_D(addr[2]),
    .Q_E(addr[1]),
    .Q_F(addr[0]),
    .Q_G(addr[10]),
    .Q_H(ba[1]),
    .Q_H_n()
);

\74595 three(
    .SER(ser3),
    .SCLK(srclk),
    .RCLK(rclk),
    .OE_n(1'b0),
    .CLR_n(1'b1),
    .VCC(1'b1),
    .GND(1'b0),
    .Q_A(dqm[0]),
    .Q_B(dqm[1]),
    .Q_C(cke),
    .Q_D(), // .Q_D(csb),
    .Q_E(rasb),
    .Q_F(casb),
    .Q_G(web),
    .Q_H(),
    .Q_H_n()
);

// logic dq_en = 0;
// logic [15:0] dq_in;
// assign dq = dq_en ? dq_in : 16'bZ;

initial begin
    $display("Starting simulation");


#0ns;  ser1 <= 0;  ser2 <= 0;  ser3 <= 0;  rclk <= 1;  clk <= 1;
#19ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  ser3 <= 1;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser3 <= 0;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  rclk <= 0;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  rclk <= 1;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser2 <= 1;  ser3 <= 1;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  ser2 <= 0;  ser3 <= 0;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  ser3 <= 1;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  ser3 <= 0;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser3 <= 1;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  rclk <= 0;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  rclk <= 1;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  ser3 <= 1;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  ser3 <= 0;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  ser3 <= 1;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  ser3 <= 0;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  rclk <= 0;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  rclk <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser3 <= 0;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser3 <= 1;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  rclk <= 0;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  rclk <= 1;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser2 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser2 <= 0;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser3 <= 1;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  rclk <= 0;  clk <= 0;
#59ns;  clk <= 1;
#69ns;  rclk <= 1;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  ser3 <= 1;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser3 <= 0;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  ser3 <= 0;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  rclk <= 0;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  rclk <= 1;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  rclk <= 0;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  ser1 <= 1;  rclk <= 1;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser1 <= 0;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser1 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  ser1 <= 0;  ser3 <= 1;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser3 <= 0;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser1 <= 1;  rclk <= 0;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser1 <= 0;  rclk <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#69ns;  ser3 <= 1;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  ser3 <= 0;  clk <= 0;
#60ns;  clk <= 1;
#60ns;  rclk <= 0;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  rclk <= 1;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  ser3 <= 1;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  ser3 <= 0;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser3 <= 1;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser3 <= 0;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  rclk <= 0;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  rclk <= 1;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  ser3 <= 1;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  ser3 <= 0;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  ser3 <= 1;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  ser3 <= 0;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  rclk <= 0;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  rclk <= 1;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser3 <= 1;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#69ns;  rclk <= 0;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  rclk <= 1;  clk <= 0;
#60ns;  clk <= 1;
#60ns;  ser2 <= 1;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser2 <= 0;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  ser3 <= 1;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  ser3 <= 0;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  ser3 <= 1;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  ser3 <= 0;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  rclk <= 0;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  rclk <= 1;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  ser3 <= 1;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser3 <= 0;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser3 <= 1;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  ser3 <= 0;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  rclk <= 0;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  rclk <= 1;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser3 <= 1;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  ser3 <= 0;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  ser3 <= 1;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser3 <= 0;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  rclk <= 0;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  rclk <= 1;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#60ns;  ser3 <= 1;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  ser3 <= 0;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  rclk <= 0;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  rclk <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser2 <= 1;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser2 <= 0;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  ser3 <= 1;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser3 <= 0;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#69ns;  rclk <= 0;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  rclk <= 1;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser3 <= 1;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  ser3 <= 1;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  ser3 <= 0;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  rclk <= 0;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  rclk <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  rclk <= 0;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  rclk <= 1;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser2 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#69ns;  ser2 <= 0;  ser3 <= 1;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  ser3 <= 0;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser3 <= 1;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  ser3 <= 0;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  rclk <= 0;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#9ns;  rclk <= 1;
#59ns;  clk <= 1;
#59ns;  ser3 <= 1;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser3 <= 0;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#10ns;  ser3 <= 1;
#59ns;  clk <= 1;
#59ns;  ser3 <= 0;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  rclk <= 0;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  rclk <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  rclk <= 0;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  ser1 <= 1;  rclk <= 1;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser1 <= 0;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#9ns;  ser1 <= 1;
#60ns;  clk <= 1;
#59ns;  ser1 <= 0;  ser3 <= 1;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser3 <= 0;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser1 <= 1;  rclk <= 0;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser1 <= 0;  rclk <= 1;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#9ns;  ser3 <= 1;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#69ns;  ser3 <= 1;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  rclk <= 0;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  rclk <= 1;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser3 <= 1;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  rclk <= 0;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#9ns;  rclk <= 1;
#60ns;  clk <= 1;
#59ns;  ser3 <= 1;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#9ns;  ser3 <= 1;
#59ns;  clk <= 1;
#60ns;  ser3 <= 0;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  rclk <= 0;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  rclk <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#60ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#70ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#60ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#60ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#60ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#70ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#70ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#60ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#60ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#70ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#9ns;  ser3 <= 1;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser3 <= 0;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  rclk <= 0;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  rclk <= 1;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser2 <= 1;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  ser2 <= 0;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#10ns;  ser3 <= 1;
#60ns;  clk <= 1;
#59ns;  ser3 <= 0;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser3 <= 1;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser3 <= 0;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  rclk <= 0;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#10ns;  rclk <= 1;
#59ns;  clk <= 1;
#59ns;  ser3 <= 1;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  ser3 <= 0;  clk <= 0;
#60ns;  clk <= 1;
#60ns;  clk <= 0;
#10ns;  ser3 <= 1;
#59ns;  clk <= 1;
#60ns;  ser3 <= 0;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  rclk <= 0;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  rclk <= 1;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  ser3 <= 1;  clk <= 0;
#60ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser3 <= 0;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#69ns;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  rclk <= 0;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  rclk <= 1;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#60ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#70ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#60ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#60ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#70ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#70ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#60ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#60ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#70ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#60ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  ser3 <= 0;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  rclk <= 0;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  rclk <= 1;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser2 <= 1;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#69ns;  ser2 <= 0;  ser3 <= 0;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  ser3 <= 1;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#9ns;  ser3 <= 0;
#59ns;  clk <= 1;
#60ns;  ser3 <= 1;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  ser3 <= 0;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  rclk <= 0;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  rclk <= 1;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#10ns;  ser3 <= 1;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#69ns;  ser3 <= 1;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#9ns;  ser3 <= 0;
#60ns;  clk <= 1;
#59ns;  rclk <= 0;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  rclk <= 1;  clk <= 0;
#59ns;  clk <= 1;
#69ns;  ser3 <= 1;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  ser3 <= 0;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser3 <= 1;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  rclk <= 0;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#9ns;  rclk <= 1;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser2 <= 1;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser2 <= 0;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#10ns;  ser3 <= 1;
#59ns;  clk <= 1;
#59ns;  ser3 <= 0;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  rclk <= 0;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  rclk <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#10ns;  ser3 <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#69ns;  ser3 <= 0;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  rclk <= 0;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  rclk <= 1;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#69ns;  ser3 <= 0;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  ser3 <= 1;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser3 <= 0;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  rclk <= 0;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser1 <= 1;  rclk <= 1;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  ser1 <= 0;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser1 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser1 <= 0;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#10ns;  ser3 <= 0;
#59ns;  clk <= 1;
#59ns;  ser1 <= 1;  rclk <= 0;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser1 <= 0;  rclk <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser3 <= 0;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  rclk <= 0;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  rclk <= 1;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser3 <= 1;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#9ns;  ser3 <= 1;
#59ns;  clk <= 1;
#60ns;  ser3 <= 0;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  rclk <= 0;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  rclk <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  rclk <= 0;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  rclk <= 1;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  ser3 <= 1;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser3 <= 0;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  ser3 <= 1;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  ser3 <= 0;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  rclk <= 0;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  rclk <= 1;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser2 <= 1;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  ser2 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#10ns;  ser3 <= 0;
#59ns;  clk <= 1;
#60ns;  ser3 <= 1;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  rclk <= 0;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  rclk <= 1;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  ser3 <= 1;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  ser3 <= 0;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  rclk <= 0;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  rclk <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser3 <= 0;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#69ns;  rclk <= 0;  clk <= 0;
#60ns;  clk <= 1;
#60ns;  rclk <= 1;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser3 <= 1;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  ser3 <= 0;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser3 <= 1;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser3 <= 0;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  rclk <= 0;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  rclk <= 1;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  ser2 <= 1;  ser3 <= 1;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser2 <= 0;  ser3 <= 0;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  ser3 <= 0;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  rclk <= 0;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  rclk <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser3 <= 0;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  rclk <= 0;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  rclk <= 1;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser3 <= 1;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#69ns;  ser3 <= 0;  clk <= 0;
#60ns;  clk <= 1;
#60ns;  ser3 <= 1;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser3 <= 0;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  rclk <= 0;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  rclk <= 1;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  ser2 <= 1;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser2 <= 0;  ser3 <= 1;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  ser3 <= 0;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  rclk <= 0;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  rclk <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  rclk <= 0;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  rclk <= 1;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser3 <= 1;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  ser3 <= 0;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  ser3 <= 1;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser3 <= 0;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  rclk <= 0;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser1 <= 1;  rclk <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser1 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser1 <= 1;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  ser1 <= 0;  ser3 <= 1;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  ser3 <= 0;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  ser1 <= 1;  rclk <= 0;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser1 <= 0;  rclk <= 1;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  ser3 <= 0;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser3 <= 1;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser3 <= 0;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  rclk <= 0;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  rclk <= 1;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  ser3 <= 1;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser3 <= 0;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  ser3 <= 0;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  rclk <= 0;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  rclk <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser3 <= 0;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  ser3 <= 1;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  ser3 <= 0;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  rclk <= 0;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  rclk <= 1;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#69ns;  clk <= 1;
#60ns;  clk <= 0;
#59ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#70ns;  clk <= 0;
#59ns;  clk <= 1;
#59ns;  ser3 <= 1;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  clk <= 0;
#70ns;  clk <= 1;
#59ns;  ser3 <= 0;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  clk <= 0;
#60ns;  clk <= 1;
#69ns;  ser3 <= 1;  clk <= 0;
#60ns;  clk <= 1;

end
endmodule