`timescale 1ns / 1ps

module test_sdram;

/*
module MT48LC8M16A2 (dq, addr, ba, clk, cke, csb, rasb, casb, web, dqm);

    parameter addr_bits =      13;
    parameter data_bits =      16;
    parameter col_bits  =       9;
    parameter mem_sizes = 2097151;                                  // 2 Meg
 
    inout     [data_bits - 1 : 0] dq;
    input     [addr_bits - 1 : 0] addr;
    input                 [1 : 0] ba;
    input                         clk;
    input                         cke;
    input                         csb;
    input                         rasb;
    input                         casb;
    input                         web;
    input                 [1 : 0] dqm;
*/

wire [15:0] dq;
logic [12:0] addr;
logic [1:0] ba;
logic clk;
logic cke;
logic csb;
logic rasb;
logic casb;
logic web;
logic [1:0] dqm;

logic srclk, rclk, ser1, ser2, ser3;

IS42VM16400K
// MT48LC8M16A2 
sdram(
    .dq(dq),
    .addr(addr),
    .ba(ba),
    .clk(clk),
    .cke(cke),
    .csb(csb),
    .rasb(rasb),
    .casb(casb),
    .web(web),
    .dqm(dqm)
);

\74595 one(
    .SER(ser1),
    .SCLK(srclk),
    .RCLK(rclk),
    .OE_n(0),
    .CLR_n(1),
    .VCC(1),
    .GND(0),
    .Q_A(addr[4]),
    .Q_B(addr[12]),
    .Q_C(addr[11]),
    .Q_D(addr[9]),
    .Q_E(addr[8]),
    .Q_F(addr[7]),
    .Q_G(addr[6]),
    .Q_H(addr[5]),
    .Q_H_n()
);

\74595 two(
    .SER(ser2),
    .SCLK(srclk),
    .RCLK(rclk),
    .OE_n(0),
    .CLR_n(1),
    .VCC(1),
    .GND(0),
    .Q_A(ba[0]),
    .Q_B(),
    .Q_C(addr[3]),
    .Q_D(addr[2]),
    .Q_E(addr[1]),
    .Q_F(addr[0]),
    .Q_G(addr[10]),
    .Q_H(ba[1]),
    .Q_H_n()
);

\74595 three(
    .SER(ser3),
    .SCLK(srclk),
    .RCLK(rclk),
    .OE_n(0),
    .CLR_n(1),
    .VCC(1),
    .GND(0),
    .Q_A(dqm[0]),
    .Q_B(dqm[1]),
    .Q_C(cke),
    .Q_D(csb),
    .Q_E(rasb),
    .Q_F(casb),
    .Q_G(web),
    .Q_H(),
    .Q_H_n()
);

// logic dq_en = 0;
// logic [15:0] dq_in;
// assign dq = dq_en ? dq_in : 16'bZ;

initial begin
    $display("Starting simulation");

#0.000ns;  ser1 <= 0;  ser2 <= 0;  ser3 <= 0;  rclk <= 0;  srclk <= 0;  clk <= 0;
#3774.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#48.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  rclk <= 1;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#8.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  rclk <= 0;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  ser3 <= 0;  rclk <= 1;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  ser2 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  ser2 <= 0;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;  clk <= 1;
#8.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  srclk <= 0;
#2.000ns;  ser3 <= 1;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#8.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser1 <= 1;  rclk <= 1;  srclk <= 0;  clk <= 0;
#8.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  ser1 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser2 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser1 <= 1;  ser2 <= 0;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#2.000ns;  ser1 <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#8.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;  clk <= 1;
#8.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#12.000ns;  rclk <= 0;
#38.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  rclk <= 1;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#8.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#2.000ns;  ser3 <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#8.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  ser2 <= 1;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  ser2 <= 0;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#8.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;  clk <= 1;
#8.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#10.000ns;  rclk <= 0;
#42.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  rclk <= 1;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#2.000ns;  ser3 <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#8.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#8.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  ser2 <= 1;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser2 <= 0;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#8.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  rclk <= 0;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  rclk <= 1;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#8.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;  clk <= 1;
#8.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  ser2 <= 1;  ser3 <= 1;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  ser2 <= 0;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  ser3 <= 0;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#8.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  rclk <= 0;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  rclk <= 1;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#8.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#8.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  ser2 <= 1;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser2 <= 0;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#8.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  rclk <= 0;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  rclk <= 1;  clk <= 0;
#8.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#8.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  ser2 <= 1;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  ser2 <= 0;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;  clk <= 1;
#8.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  ser3 <= 1;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#2.000ns;  rclk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  rclk <= 1;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;  clk <= 1;
#8.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  ser3 <= 1;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#8.000ns;  ser2 <= 1;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser2 <= 0;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#8.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  rclk <= 0;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  rclk <= 1;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#8.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#8.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  ser2 <= 1;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#2.000ns;  ser2 <= 0;  ser3 <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#8.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;  clk <= 1;
#8.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#2.000ns;  rclk <= 0;
#50.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  rclk <= 1;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#8.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;  clk <= 1;
#8.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  ser2 <= 1;  ser3 <= 1;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  ser2 <= 0;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  ser3 <= 0;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#8.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#6.000ns;  rclk <= 0;
#44.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  rclk <= 1;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#8.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#8.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  ser2 <= 1;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser2 <= 0;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#8.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  rclk <= 0;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  rclk <= 1;  clk <= 0;
#8.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#8.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  ser2 <= 1;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  ser2 <= 0;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;  clk <= 1;
#8.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  ser3 <= 1;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#2.000ns;  rclk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  rclk <= 1;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;  clk <= 1;
#8.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  ser3 <= 1;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#8.000ns;  ser2 <= 1;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser2 <= 0;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#8.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  rclk <= 0;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  rclk <= 1;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#8.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#8.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  ser2 <= 1;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#2.000ns;  ser2 <= 0;  ser3 <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#8.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;  clk <= 1;
#8.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#50.000ns;  clk <= 1;
#52.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#2.000ns;  rclk <= 0;
#50.000ns;  clk <= 1;
#50.000ns;  clk <= 0;
#52.000ns;  clk <= 1;
#52.000ns;  rclk <= 1;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;  clk <= 1;
#6.000ns;  srclk <= 1;
#8.000ns;  ser3 <= 1;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 0;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#8.000ns;  srclk <= 1;
#6.000ns;  rclk <= 1;  srclk <= 0;  clk <= 0;
#6.000ns;  rclk <= 0;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#8.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
#6.000ns;  srclk <= 1;
#6.000ns;  ser3 <= 1;  srclk <= 0;  clk <= 1;
#8.000ns;  srclk <= 1;
#6.000ns;  srclk <= 0;
end
endmodule